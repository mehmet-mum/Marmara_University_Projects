module control(in,regdest,alusrc,memtoreg,regwrite,memread,memwrite,branch,aluop1,aluop2,jump,b_new,flag,link,addr_from_mem);
input [5:0] in;
output regdest,alusrc,memtoreg,regwrite,memread,memwrite,branch,aluop1,aluop2,jump,b_new,link,addr_from_mem;
output [1:0] flag;
wire rformat,lw,sw,beq,bmn,bz,jalm,jump_ins;
assign rformat=~|in;
assign lw=in[5]& (~in[4])&(~in[3])&(~in[2])&in[1]&in[0];
assign sw=in[5]& (~in[4])&in[3]&(~in[2])&in[1]&in[0];
assign beq=~in[5]& (~in[4])&(~in[3])&in[2]&(~in[1])&(~in[0]);
assign bmn=~in[5]& in[4] & (~in[3]) & in[2] & (~in[1]) & in[0];
assign bz=~in[5]& in[4] & in[3] & (~in[2]) & (~in[1]) & (~in[0]);
assign jalm=~in[5]& in[4] & (~in[3])& (~in[2]) & in[1] & in[0];
assign jump_ins=(~in[5])&(~in[4])&(~in[3])&(~in[2])&(in[1])&(~in[0]);
assign regdest=rformat;
assign alusrc=lw|sw|bmn|jalm;
assign memtoreg=lw|jalm|bmn;
assign regwrite=rformat|lw|jalm;
assign memread=lw|bmn|jalm;
assign memwrite=sw;
assign branch=beq|jalm|bmn;
assign aluop1=rformat;
assign aluop2=beq;
assign b_new=rformat|bmn|bz|jalm;
assign flag[1]= bmn;
assign flag[0]=jalm;
assign link=jalm;
assign jump=jump_ins|bz;
assign addr_from_mem=jalm|rformat|bmn;
endmodule
